module AND_GATE(C, A,B);
	input A,B;
	output C;
	assign C = A & B;
endmodule